`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2019/03/09 19:51:29
// Design Name: 
// Module Name: test_frequency_divider_about_1hz
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module test_frequency_divider_about_1hz;
    reg [26:0] q;
    wire clk, rst;
    initial begin
        clk = 1'b0;
    end
endmodule
